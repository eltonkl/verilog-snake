module Debouncer(
    input wire 	Clock,
    input wire  Signal,
    output wire Pressed
    );


endmodule
