`include "Constants.v"

module Snake(
    input wire          ButtonLeft,
    input wire          ButtonRight,
    input wire          ButtonUp,
    input wire          ButtonDown,
    input wire          ButtonCenter,
    output wire [0:2]   VGARed,
    output wire [0:2]   VGAGreen,
    output wire [0:1]   VGABlue,
    output wire         VGAHSync,
    output wire         VGAVSync
    );


endmodule
