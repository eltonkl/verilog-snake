`include "Constants.vh"

module VGAController(
    output reg [0:2]    Red,
    output reg [0:2]    Green,
    output reg [0:1]    Blue,
    output              HSync,
    output              VSync
    );


endmodule
